module LED(i, j);

input i;
output j;

assign j = i;

endmodule



